library ieee;
use ieee.std_logic_1164.all;


entity full_adder is
port(
	x, y, cin : in std_logic;
	s, cout : out std_logic
	);
	
	
end full_adder;

architecture rtl of full_adder is
begin

	s <= x xor y xor cin;
	cout <= (x and y) or (x and cin) or (y and cin);
	
	
end rtl;